module template();

endmodule
