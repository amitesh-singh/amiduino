module led(output led1, output led2, output led3, output led4);
//input s1; // Location: PIN_88, I/O Standard: 3.3-V LVTTL, Current Strength: 8mA
//input s2; // Location: PIN_89, I/O Standard: 3.3-V LVTTL, Current Strength: 8mA
	//output led1; // Location: PIN_87, I/O Standard: 3.3-V LVTTL, Current Strength: 8mA
	assign led1 = 0; //this will switch on the led1
	assign led2 = 0; //this will switch on the led2
	assign led3 = 0; //this will switch on the led3
	assign led4 = 0; //this will switch on the led4
endmodule